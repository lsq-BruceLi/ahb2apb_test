woshui jdkfjd



lidada



2023年 10月 30日 星期一 16:17:09 CST
