hfah





2023年 10月 30日 星期一 16:19:47 CST
